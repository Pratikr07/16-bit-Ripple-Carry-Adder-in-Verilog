module adder16bit(x,y,z,sign,zero,carry,parity,overflow);

   input [15:0]x,y;
   output [15:0]z;
   output sign,zero,carry,parity,overflow;
   wire [3:1]c;

   assign sign= z[15];
   assign zero= ~|z;
   assign parity= ~^z;
   assign overflow= (x[15] & y[15] & ~z[15]) | (~x[15] & ~y[15] & z[15]);

   adder4bit A0 (z[3:0],c[1],x[3:0],y[3:0],1'b0);
   adder4bit A1 (z[7:4],c[2],x[7:4],y[7:4],c[1]);
   adder4bit A2 (z[11:8],c[3],x[11:8],y[11:8],c[2]);
   adder4bit A3 (z[15:12],carry,x[15:12],y[15:12],c[3]);

endmodule